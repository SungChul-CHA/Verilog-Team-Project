`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// ne u (.a(), .b(), .o());
// Not Equal -> 1 Equal -> 0
// Maker : CHA
//
//////////////////////////////////////////////////////////////////////////////////


module ne(
    input a,
    input b,
    output reg o
    );
    
    always @ (a or b) begin
        if (a!=b) o = 1;
        else o = 0;
    end
    
endmodule
