`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// ge u (.a(), .b(), .o());
// a >= b -> 1
// Maker : CHA
//
//////////////////////////////////////////////////////////////////////////////////


module ge(
    input a,
    input b,
    output reg o
    );
    
    always @ (a or b) begin
        if (a >= b) o = 1;
        else o = 0;
    end
    
endmodule
