`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// eq u (.a(), .b(), .o());
// Equal -> 1 Not Equal -> 0
// Maker : CHA
//
//////////////////////////////////////////////////////////////////////////////////


module eq(
    input a,
    input b,
    output reg o
    );
    
    always @ (a or b) begin
        if (a == b) o = 1;
        else o = 0;
    end
    
endmodule
